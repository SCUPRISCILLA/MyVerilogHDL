module my3_8code(a, b, c, l);
input a, b, c;
output reg[7:0] l;

always@(*)
begin
case({c, b, a})
3'b000: l <= 8'b0000_0001;
3'b001: l <= 8'b0000_0010;
3'b010: l <= 8'b0000_0100;
3'b011: l <= 8'b0000_1000;
3'b100: l <= 8'b0001_0000;
3'b101: l <= 8'b0010_0000;
3'b110: l <= 8'b0100_0000;
3'b111: l <= 8'b1000_0000;
endcase
end
endmodule